----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:55:17 03/26/2018 
-- Design Name: 
-- Module Name:    adder4 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity adder4 is
    Port ( i_a : in  STD_LOGIC_VECTOR (3 downto 0);
           i_b : in  STD_LOGIC_VECTOR (3 downto 0);
           i_c : in  STD_LOGIC;
           o_out : out  STD_LOGIC_VECTOR (3 downto 0);
           o_c : out  STD_LOGIC);
end adder4;

architecture Behavioral of adder4 is

begin


end Behavioral;

